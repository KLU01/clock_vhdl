library verilog;
use verilog.vl_types.all;
entity mod6_vlg_vec_tst is
end mod6_vlg_vec_tst;
