library verilog;
use verilog.vl_types.all;
entity BCD_Counter3_vlg_vec_tst is
end BCD_Counter3_vlg_vec_tst;
